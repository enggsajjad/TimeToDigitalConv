library verilog;
use verilog.vl_types.all;
entity top_drom_tf is
end top_drom_tf;
