library verilog;
use verilog.vl_types.all;
entity testcounter_tf_v_tf is
end testcounter_tf_v_tf;
