library verilog;
use verilog.vl_types.all;
entity cu_hmi_tf is
end cu_hmi_tf;
