library verilog;
use verilog.vl_types.all;
entity chrono48_start_tf is
end chrono48_start_tf;
