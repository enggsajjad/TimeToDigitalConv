library verilog;
use verilog.vl_types.all;
entity ir_decoder_tf is
end ir_decoder_tf;
